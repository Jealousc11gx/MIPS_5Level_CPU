//write back
//`include "define.v"

//module wb (
//***************
//);
//***************    
//endmodule